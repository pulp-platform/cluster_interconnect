`ifndef MUT_IMPL
  `define MUT_IMPL 1
 `endif
`ifndef NUM_MASTER
  `define NUM_MASTER 64
 `endif
`ifndef BANK_FACT
  `define BANK_FACT 1
 `endif
`ifndef DATA_WIDTH
  `define DATA_WIDTH 32
`endif
`ifndef MEM_ADDR_BITS
  `define MEM_ADDR_BITS 12
`endif
`ifndef PAR_STAGES
  `define PAR_STAGES 1
`endif
`ifndef TEST_CYCLES
  `define TEST_CYCLES 2000
`endif
